module dmem(
    input clk,
    input MemRW,
    input [31:0] addr,
    input [31:0] dataW,
    input [3:0] MemWriteMask,
    output [31:0] dataR
);


endmodule